
import MicroSD::*;
import Conv2D::*;
import BatchPool::*;
import FRAM::*;



interface WildfireIfc;

endinterface

module mkWildfire(WildfireIfc);







endmodule
